`ifndef PRIMITIVE_TYPES_SVH
`define PRIMITIVE_TYPES_SVH
package primitive_types;
    typedef logic [7:0] node_id_t;
    typedef logic [7:0] packet_id_t;
    typedef logic [7:0] flit_num_t;
endpackage
`endif
