module flit_buffer();
endmodule
