module noc();
endmodule
