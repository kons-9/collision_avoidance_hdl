module packet_transfer_buffer();
  // MUST TODO
  // 完了したパケットの送信を担当する
endmodule
