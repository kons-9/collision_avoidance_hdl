module ack_controller();
endmodule
