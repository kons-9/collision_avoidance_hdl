/// 通常のフリットの場合、ACKを生成するモジュール
module make_ack_comb(
    input types::flit_t flit_in,
    input logic flit_in_vld,

    output types::flit_t flit_out,
    output logic flit_out_vld
);
// TODO

endmodule
