/// 通常のフリットの場合、ACKを生成するモジュール
module make_ack_comb(
    input types::flit_t flit_in,

    output types::flit_t flit_out
);
// MUST TODO

endmodule
