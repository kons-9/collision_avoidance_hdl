module combine_flit (
    input logic clk,
    input logic rst_n,

    output types::flit_t flit_out,
    output logic  flit_out_vld
);
  // TODO
endmodule
