module uart_rx (
    input  logic  uart_clk,
    input  logic  rst_n,
    input  logic  uart_rx,
    output flit_t flit_out,
    output logic  flit_out_vld
);
endmodule
