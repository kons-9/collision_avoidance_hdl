module receive_controller();
endmodule
