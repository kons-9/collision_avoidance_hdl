`include "types.svh"
