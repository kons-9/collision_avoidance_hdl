/// 受信したデータのヘッダーを見て、適切な信号処理を行う
module control_received_flit ();
  // TODO: 現在の実装はack待ちをブロッキングで行う予定
  // 将来的にはack待ちbufferを作成する
endmodule
