/// ack, sendの優先度でflitを取り出す
module pop_flit ();
  // TODO
endmodule
