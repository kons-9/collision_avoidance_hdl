module uart_tx (
    input  logic  uart_clk,
    input  logic  rst_n,
    input  logic  flit_in_vld,
    input  flit_t flit_in,
    output logic  flit_in_rdy
);
endmodule
