module buffer_update(
  input buffer_t rx_buffer,

  

);

endmodule
